<ion-menu [content]="content">
    <ion-header>
        <ion-toolbar>
            <ion-title>Menu</ion-title>
        </ion-toolbar>
    </ion-header>

    <ion-content>
        <ion-list>
            <button ion-item (click)="onHomeButtonClicked()">
                <ion-icon name="home_" item-start></ion-icon>
                <ion-label>Home</ion-label>
            </button>
            <button *ngIf="this.localStorageProvider.isUserRegistered()" ion-item (click)="onFavoritesButtonClicked()">
                <ion-icon name="favorite_" item-start></ion-icon>
                <ion-label>Favorites</ion-label>
            </button>
            <button *ngIf="this.localStorageProvider.isUserRegistered()" ion-item (click)="onWalletsButtonClicked()">
                <ion-icon name="wallet_" item-start></ion-icon>
                <ion-label>Wallets</ion-label>
            </button>
            <button *ngIf="this.localStorageProvider.isUserRegistered()" ion-item (click)="onAlertsButtonClicked()">
                <ion-icon name="alert_" item-start></ion-icon>
                <ion-label>Alerts</ion-label>
            </button>
            <button *ngIf="this.localStorageProvider.isUserRegistered()" ion-item (click)="onSettingsButtonClicked()">
                <ion-icon name="setting_" item-start></ion-icon>
                <ion-label>Settings</ion-label>
            </button>
            <button *ngIf="!this.localStorageProvider.isUserRegistered()" ion-item (click)="onSubscribeButtonClicked()">
                <ion-icon name="subscribe_" item-start></ion-icon>
                <ion-label>Subscribe</ion-label>
            </button>
            <button *ngIf="!this.localStorageProvider.isUserRegistered()" ion-item (click)="onLogInButtonClicked()">
                <ion-icon name="log-in_" item-start></ion-icon>
                <ion-label>Log in</ion-label>
            </button>
        </ion-list>
    </ion-content>
</ion-menu>

<ion-nav #content [root]="rootPage"></ion-nav>